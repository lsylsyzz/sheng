module add3(a,
b,
c,
cout);

input [2:0] a,b;
input cout;
output [2:0]c;
///assign c=a+b;
//assign cout = (a[2]==b[2])&&(c[2] != b[2])?1:0;

endmodule
