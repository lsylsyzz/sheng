module top_module( 
    input [99:0] a, b,
    input sel,
    output [99:0] out );

   wire sel ;
   // assign out = sel ? b : a;
endmodule

